

library ieee;
library work;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
use work.fft_types.all;

-- delay is 5 cycles

entity windowMultiply1024_64 is
	generic(dataBits, outBits: integer := 18);
	port(clk: in std_logic;
			din: in complex;
			index: in unsigned(10-1 downto 0);
			dout: out complex
			);
end entity;
architecture a of windowMultiply1024_64 is
	constant romDepthOrder: integer := 10;
	constant romDepth: integer := 2**romDepthOrder;
	constant romWidth: integer := 18;
	--ram
	type ram1t is array(0 to romDepth-1) of
		std_logic_vector(romWidth-1 downto 0);
	signal rom: ram1t;
	signal addr1: unsigned(romDepthOrder-1 downto 0);
	signal data0, data1, data2: std_logic_vector(romWidth-1 downto 0);
	signal coeff: signed(romWidth-1 downto 0);

	signal din1, din2, din3: complex;

	-- multiplier
	signal multOutRe, multOutIm: signed(dataBits+romWidth-1 downto 0);
	signal multOut, multOut1: complex;

	attribute keep: string;
	attribute keep of din2: signal is "true";
	attribute keep of data2: signal is "true";
begin
	-- coefficient rom
	addr1 <= index; -- when rising_edge(clk);
	data0 <= rom(to_integer(addr1));
	data1 <= data0 when rising_edge(clk);
	data2 <= data1 when rising_edge(clk);
	coeff <= signed(data2) when rising_edge(clk);

	-- delay data
	din1 <= din when rising_edge(clk);
	din2 <= din1 when rising_edge(clk);
	din3 <= din2 when rising_edge(clk);

	-- multiply
	multOutRe <= coeff * complex_re(din3, dataBits);
	multOutIm <= coeff * complex_im(din3, dataBits);

	multOut <= to_complex(multOutRe(multOutRe'left-1 downto multOutRe'left-outBits),
						multOutIm(multOutIm'left-1 downto multOutIm'left-outBits));
	multOut1 <= multOut when rising_edge(clk);
	dout <= multOut1 when rising_edge(clk);

	-- rom
	rom <= (

"000000000000000000" , "000000000000000000" , "000000000000000000" , "000000000000000000" , "111111111111111111" , "111111111111111111" , "111111111111111111" , "111111111111111111" , "111111111111111111" , "111111111111111111" ,
"111111111111111111" , "111111111111111111" , "111111111111111111" , "111111111111111111" , "111111111111111111" , "111111111111111111" , "111111111111111111" , "111111111111111111" , "111111111111111111" , "111111111111111110" ,
"111111111111111110" , "111111111111111110" , "111111111111111110" , "111111111111111110" , "111111111111111110" , "111111111111111110" , "111111111111111110" , "111111111111111110" , "111111111111111110" , "111111111111111110" ,
"111111111111111110" , "111111111111111110" , "111111111111111110" , "111111111111111110" , "111111111111111110" , "111111111111111110" , "111111111111111110" , "111111111111111110" , "111111111111111111" , "111111111111111111" ,
"111111111111111111" , "111111111111111111" , "111111111111111111" , "000000000000000000" , "000000000000000000" , "000000000000000001" , "000000000000000001" , "000000000000000001" , "000000000000000010" , "000000000000000011" ,
"000000000000000011" , "000000000000000100" , "000000000000000101" , "000000000000000101" , "000000000000000110" , "000000000000000111" , "000000000000001000" , "000000000000001001" , "000000000000001010" , "000000000000001011" ,
"000000000000001100" , "000000000000001101" , "000000000000001111" , "000000000000010000" , "000000000000010001" , "000000000000010011" , "000000000000010100" , "000000000000010110" , "000000000000010111" , "000000000000011001" ,
"000000000000011011" , "000000000000011101" , "000000000000011111" , "000000000000100000" , "000000000000100010" , "000000000000100100" , "000000000000100111" , "000000000000101001" , "000000000000101011" , "000000000000101101" ,
"000000000000101111" , "000000000000110010" , "000000000000110100" , "000000000000110110" , "000000000000111001" , "000000000000111011" , "000000000000111110" , "000000000001000000" , "000000000001000010" , "000000000001000101" ,
"000000000001000111" , "000000000001001010" , "000000000001001100" , "000000000001001110" , "000000000001010001" , "000000000001010011" , "000000000001010101" , "000000000001010111" , "000000000001011010" , "000000000001011100" ,
"000000000001011101" , "000000000001011111" , "000000000001100001" , "000000000001100011" , "000000000001100100" , "000000000001100101" , "000000000001100111" , "000000000001101000" , "000000000001101000" , "000000000001101001" ,
"000000000001101001" , "000000000001101010" , "000000000001101010" , "000000000001101001" , "000000000001101001" , "000000000001101000" , "000000000001100111" , "000000000001100110" , "000000000001100100" , "000000000001100010" ,
"000000000001100000" , "000000000001011110" , "000000000001011011" , "000000000001010111" , "000000000001010100" , "000000000001010000" , "000000000001001011" , "000000000001000110" , "000000000001000001" , "000000000000111011" ,
"000000000000110101" , "000000000000101110" , "000000000000100111" , "000000000000100000" , "000000000000011000" , "000000000000001111" , "000000000000000110" , "111111111111111100" , "111111111111110010" , "111111111111101000" ,
"111111111111011101" , "111111111111010001" , "111111111111000101" , "111111111110111001" , "111111111110101011" , "111111111110011110" , "111111111110010000" , "111111111110000001" , "111111111101110010" , "111111111101100010" ,
"111111111101010010" , "111111111101000001" , "111111111100110000" , "111111111100011110" , "111111111100001100" , "111111111011111010" , "111111111011100111" , "111111111011010011" , "111111111011000000" , "111111111010101011" ,
"111111111010010111" , "111111111010000010" , "111111111001101101" , "111111111001011000" , "111111111001000010" , "111111111000101100" , "111111111000010110" , "111111111000000000" , "111111110111101010" , "111111110111010011" ,
"111111110110111101" , "111111110110100110" , "111111110110010000" , "111111110101111010" , "111111110101100011" , "111111110101001101" , "111111110100110111" , "111111110100100010" , "111111110100001101" , "111111110011111000" ,
"111111110011100011" , "111111110011001111" , "111111110010111100" , "111111110010101001" , "111111110010010111" , "111111110010000101" , "111111110001110100" , "111111110001100100" , "111111110001010101" , "111111110001000111" ,
"111111110000111010" , "111111110000101110" , "111111110000100011" , "111111110000011001" , "111111110000010001" , "111111110000001010" , "111111110000000100" , "111111110000000000" , "111111101111111101" , "111111101111111100" ,
"111111101111111100" , "111111101111111111" , "111111110000000011" , "111111110000001000" , "111111110000010000" , "111111110000011010" , "111111110000100110" , "111111110000110100" , "111111110001000100" , "111111110001010110" ,
"111111110001101010" , "111111110010000001" , "111111110010011010" , "111111110010110110" , "111111110011010011" , "111111110011110100" , "111111110100010111" , "111111110100111100" , "111111110101100100" , "111111110110001111" ,
"111111110110111100" , "111111110111101100" , "111111111000011110" , "111111111001010100" , "111111111010001100" , "111111111011000110" , "111111111100000100" , "111111111101000100" , "111111111110000110" , "111111111111001100" ,
"000000000000010100" , "000000000001011111" , "000000000010101100" , "000000000011111100" , "000000000101001110" , "000000000110100011" , "000000000111111010" , "000000001001010100" , "000000001010110000" , "000000001100001111" ,
"000000001101101111" , "000000001111010010" , "000000010000110110" , "000000010010011101" , "000000010100000101" , "000000010101101111" , "000000010111011011" , "000000011001001000" , "000000011010110111" , "000000011100100111" ,
"000000011110011000" , "000000100000001010" , "000000100001111101" , "000000100011110000" , "000000100101100100" , "000000100111011001" , "000000101001001101" , "000000101011000010" , "000000101100110111" , "000000101110101011" ,
"000000110000011110" , "000000110010010001" , "000000110100000011" , "000000110101110100" , "000000110111100100" , "000000111001010010" , "000000111010111110" , "000000111100101000" , "000000111110010000" , "000000111111110110" ,
"000001000001011001" , "000001000010111001" , "000001000100010101" , "000001000101101111" , "000001000111000101" , "000001001000010111" , "000001001001100101" , "000001001010101110" , "000001001011110011" , "000001001100110011" ,
"000001001101101110" , "000001001110100100" , "000001001111010100" , "000001001111111111" , "000001010000100011" , "000001010001000001" , "000001010001011000" , "000001010001101001" , "000001010001110011" , "000001010001110110" ,
"000001010001110001" , "000001010001100100" , "000001010001010000" , "000001010000110100" , "000001010000001111" , "000001001111100010" , "000001001110101100" , "000001001101101110" , "000001001100100110" , "000001001011010110" ,
"000001001001111100" , "000001001000011001" , "000001000110101100" , "000001000100110110" , "000001000010110110" , "000001000000101100" , "000000111110011000" , "000000111011111010" , "000000111001010010" , "000000110110100000" ,
"000000110011100100" , "000000110000011110" , "000000101101001101" , "000000101001110011" , "000000100110001110" , "000000100010011111" , "000000011110100110" , "000000011010100011" , "000000010110010110" , "000000010001111111" ,
"000000001101011111" , "000000001000110101" , "000000000100000010" , "111111111111000110" , "111111111010000000" , "111111110100110010" , "111111101111011011" , "111111101001111100" , "111111100100010101" , "111111011110100110" ,
"111111011000110000" , "111111010010110010" , "111111001100101110" , "111111000110100011" , "111111000000010010" , "111110111001111011" , "111110110011011111" , "111110101100111110" , "111110100110011001" , "111110011111101111" ,
"111110011001000011" , "111110010010010011" , "111110001011100000" , "111110000100101100" , "111101111101110110" , "111101110111000000" , "111101110000001001" , "111101101001010010" , "111101100010011101" , "111101011011101001" ,
"111101010100110111" , "111101001110001000" , "111101000111011100" , "111101000000110101" , "111100111010010010" , "111100110011110101" , "111100101101011110" , "111100100111001111" , "111100100001000110" , "111100011011000111" ,
"111100010101010000" , "111100001111100100" , "111100001010000010" , "111100000100101011" , "111011111111100001" , "111011111010100100" , "111011110101110100" , "111011110001010011" , "111011101101000001" , "111011101001000000" ,
"111011100101001111" , "111011100001110000" , "111011011110100011" , "111011011011101001" , "111011011001000011" , "111011010110110010" , "111011010100110110" , "111011010011010000" , "111011010010000001" , "111011010001001010" ,
"111011010000101011" , "111011010000100100" , "111011010000111000" , "111011010001100110" , "111011010010101111" , "111011010100010011" , "111011010110010100" , "111011011000110010" , "111011011011101101" , "111011011111000110" ,
"111011100010111110" , "111011100111010100" , "111011101100001011" , "111011110001100001" , "111011110111011000" , "111011111101110000" , "111100000100101001" , "111100001100000100" , "111100010100000001" , "111100011100100001" ,
"111100100101100011" , "111100101111001000" , "111100111001010001" , "111101000011111100" , "111101001111001100" , "111101011010111111" , "111101100111010110" , "111101110100010000" , "111110000001101111" , "111110001111110010" ,
"111110011110011000" , "111110101101100010" , "111110111101010000" , "111111001101100010" , "111111011110010111" , "111111101111101111" , "000000000001101010" , "000000010100000111" , "000000100111000111" , "000000111010101001" ,
"000001001110101100" , "000001100011010000" , "000001111000010101" , "000010001101111010" , "000010100011111111" , "000010111010100010" , "000011010001100100" , "000011101001000011" , "000100000001000000" , "000100011001011000" ,
"000100110010001100" , "000101001011011011" , "000101100101000011" , "000101111111000100" , "000110011001011110" , "000110110100001110" , "000111001111010101" , "000111101010110000" , "001000000110100000" , "001000100010100010" ,
"001000111110110111" , "001001011011011100" , "001001111000010001" , "001010010101010100" , "001010110010100101" , "001011010000000010" , "001011101101101001" , "001100001011011010" , "001100101001010011" , "001101000111010100" ,
"001101100101011001" , "001110000011100011" , "001110100001110000" , "001110111111111111" , "001111011110001110" , "001111111100011011" , "010000011010100110" , "010000111000101100" , "010001010110101110" , "010001110100101000" ,
"010010010010011010" , "010010110000000010" , "010011001101011111" , "010011101010101111" , "010100000111110001" , "010100100100100100" , "010101000001000101" , "010101011101010101" , "010101111001010000" , "010110010100110110" ,
"010110110000000110" , "010111001010111101" , "010111100101011011" , "010111111111011111" , "011000011001000110" , "011000110010010000" , "011001001010111011" , "011001100011000110" , "011001111010101111" , "011010010001110111" ,
"011010101000011010" , "011010111110011001" , "011011010011110001" , "011011101000100010" , "011011111100101011" , "011100010000001010" , "011100100010111111" , "011100110101001000" , "011101000110100101" , "011101010111010101" ,
"011101100111010110" , "011101110110101000" , "011110000101001010" , "011110010010111011" , "011110011111111011" , "011110101100001000" , "011110110111100010" , "011111000010001001" , "011111001011111100" , "011111010100111010" ,
"011111011101000011" , "011111100100010110" , "011111101010110011" , "011111110000011010" , "011111110101001010" , "011111111001000011" , "011111111100000101" , "011111111110010000" , "011111111111100011" , "011111111111111111" ,
"011111111111100011" , "011111111110010000" , "011111111100000101" , "011111111001000011" , "011111110101001010" , "011111110000011010" , "011111101010110011" , "011111100100010110" , "011111011101000011" , "011111010100111010" ,
"011111001011111100" , "011111000010001001" , "011110110111100010" , "011110101100001000" , "011110011111111011" , "011110010010111011" , "011110000101001010" , "011101110110101000" , "011101100111010110" , "011101010111010101" ,
"011101000110100101" , "011100110101001000" , "011100100010111111" , "011100010000001010" , "011011111100101011" , "011011101000100010" , "011011010011110001" , "011010111110011001" , "011010101000011010" , "011010010001110111" ,
"011001111010101111" , "011001100011000110" , "011001001010111011" , "011000110010010000" , "011000011001000110" , "010111111111011111" , "010111100101011011" , "010111001010111101" , "010110110000000110" , "010110010100110110" ,
"010101111001010000" , "010101011101010101" , "010101000001000101" , "010100100100100100" , "010100000111110001" , "010011101010101111" , "010011001101011111" , "010010110000000010" , "010010010010011010" , "010001110100101000" ,
"010001010110101110" , "010000111000101100" , "010000011010100110" , "001111111100011011" , "001111011110001110" , "001110111111111111" , "001110100001110000" , "001110000011100011" , "001101100101011001" , "001101000111010100" ,
"001100101001010011" , "001100001011011010" , "001011101101101001" , "001011010000000010" , "001010110010100101" , "001010010101010100" , "001001111000010001" , "001001011011011100" , "001000111110110111" , "001000100010100010" ,
"001000000110100000" , "000111101010110000" , "000111001111010101" , "000110110100001110" , "000110011001011110" , "000101111111000100" , "000101100101000011" , "000101001011011011" , "000100110010001100" , "000100011001011000" ,
"000100000001000000" , "000011101001000011" , "000011010001100100" , "000010111010100010" , "000010100011111111" , "000010001101111010" , "000001111000010101" , "000001100011010000" , "000001001110101100" , "000000111010101001" ,
"000000100111000111" , "000000010100000111" , "000000000001101010" , "111111101111101111" , "111111011110010111" , "111111001101100010" , "111110111101010000" , "111110101101100010" , "111110011110011000" , "111110001111110010" ,
"111110000001101111" , "111101110100010000" , "111101100111010110" , "111101011010111111" , "111101001111001100" , "111101000011111100" , "111100111001010001" , "111100101111001000" , "111100100101100011" , "111100011100100001" ,
"111100010100000001" , "111100001100000100" , "111100000100101001" , "111011111101110000" , "111011110111011000" , "111011110001100001" , "111011101100001011" , "111011100111010100" , "111011100010111110" , "111011011111000110" ,
"111011011011101101" , "111011011000110010" , "111011010110010100" , "111011010100010011" , "111011010010101111" , "111011010001100110" , "111011010000111000" , "111011010000100100" , "111011010000101011" , "111011010001001010" ,
"111011010010000001" , "111011010011010000" , "111011010100110110" , "111011010110110010" , "111011011001000011" , "111011011011101001" , "111011011110100011" , "111011100001110000" , "111011100101001111" , "111011101001000000" ,
"111011101101000001" , "111011110001010011" , "111011110101110100" , "111011111010100100" , "111011111111100001" , "111100000100101011" , "111100001010000010" , "111100001111100100" , "111100010101010000" , "111100011011000111" ,
"111100100001000110" , "111100100111001111" , "111100101101011110" , "111100110011110101" , "111100111010010010" , "111101000000110101" , "111101000111011100" , "111101001110001000" , "111101010100110111" , "111101011011101001" ,
"111101100010011101" , "111101101001010010" , "111101110000001001" , "111101110111000000" , "111101111101110110" , "111110000100101100" , "111110001011100000" , "111110010010010011" , "111110011001000011" , "111110011111101111" ,
"111110100110011001" , "111110101100111110" , "111110110011011111" , "111110111001111011" , "111111000000010010" , "111111000110100011" , "111111001100101110" , "111111010010110010" , "111111011000110000" , "111111011110100110" ,
"111111100100010101" , "111111101001111100" , "111111101111011011" , "111111110100110010" , "111111111010000000" , "111111111111000110" , "000000000100000010" , "000000001000110101" , "000000001101011111" , "000000010001111111" ,
"000000010110010110" , "000000011010100011" , "000000011110100110" , "000000100010011111" , "000000100110001110" , "000000101001110011" , "000000101101001101" , "000000110000011110" , "000000110011100100" , "000000110110100000" ,
"000000111001010010" , "000000111011111010" , "000000111110011000" , "000001000000101100" , "000001000010110110" , "000001000100110110" , "000001000110101100" , "000001001000011001" , "000001001001111100" , "000001001011010110" ,
"000001001100100110" , "000001001101101110" , "000001001110101100" , "000001001111100010" , "000001010000001111" , "000001010000110100" , "000001010001010000" , "000001010001100100" , "000001010001110001" , "000001010001110110" ,
"000001010001110011" , "000001010001101001" , "000001010001011000" , "000001010001000001" , "000001010000100011" , "000001001111111111" , "000001001111010100" , "000001001110100100" , "000001001101101110" , "000001001100110011" ,
"000001001011110011" , "000001001010101110" , "000001001001100101" , "000001001000010111" , "000001000111000101" , "000001000101101111" , "000001000100010101" , "000001000010111001" , "000001000001011001" , "000000111111110110" ,
"000000111110010000" , "000000111100101000" , "000000111010111110" , "000000111001010010" , "000000110111100100" , "000000110101110100" , "000000110100000011" , "000000110010010001" , "000000110000011110" , "000000101110101011" ,
"000000101100110111" , "000000101011000010" , "000000101001001101" , "000000100111011001" , "000000100101100100" , "000000100011110000" , "000000100001111101" , "000000100000001010" , "000000011110011000" , "000000011100100111" ,
"000000011010110111" , "000000011001001000" , "000000010111011011" , "000000010101101111" , "000000010100000101" , "000000010010011101" , "000000010000110110" , "000000001111010010" , "000000001101101111" , "000000001100001111" ,
"000000001010110000" , "000000001001010100" , "000000000111111010" , "000000000110100011" , "000000000101001110" , "000000000011111100" , "000000000010101100" , "000000000001011111" , "000000000000010100" , "111111111111001100" ,
"111111111110000110" , "111111111101000100" , "111111111100000100" , "111111111011000110" , "111111111010001100" , "111111111001010100" , "111111111000011110" , "111111110111101100" , "111111110110111100" , "111111110110001111" ,
"111111110101100100" , "111111110100111100" , "111111110100010111" , "111111110011110100" , "111111110011010011" , "111111110010110110" , "111111110010011010" , "111111110010000001" , "111111110001101010" , "111111110001010110" ,
"111111110001000100" , "111111110000110100" , "111111110000100110" , "111111110000011010" , "111111110000010000" , "111111110000001000" , "111111110000000011" , "111111101111111111" , "111111101111111100" , "111111101111111100" ,
"111111101111111101" , "111111110000000000" , "111111110000000100" , "111111110000001010" , "111111110000010001" , "111111110000011001" , "111111110000100011" , "111111110000101110" , "111111110000111010" , "111111110001000111" ,
"111111110001010101" , "111111110001100100" , "111111110001110100" , "111111110010000101" , "111111110010010111" , "111111110010101001" , "111111110010111100" , "111111110011001111" , "111111110011100011" , "111111110011111000" ,
"111111110100001101" , "111111110100100010" , "111111110100110111" , "111111110101001101" , "111111110101100011" , "111111110101111010" , "111111110110010000" , "111111110110100110" , "111111110110111101" , "111111110111010011" ,
"111111110111101010" , "111111111000000000" , "111111111000010110" , "111111111000101100" , "111111111001000010" , "111111111001011000" , "111111111001101101" , "111111111010000010" , "111111111010010111" , "111111111010101011" ,
"111111111011000000" , "111111111011010011" , "111111111011100111" , "111111111011111010" , "111111111100001100" , "111111111100011110" , "111111111100110000" , "111111111101000001" , "111111111101010010" , "111111111101100010" ,
"111111111101110010" , "111111111110000001" , "111111111110010000" , "111111111110011110" , "111111111110101011" , "111111111110111001" , "111111111111000101" , "111111111111010001" , "111111111111011101" , "111111111111101000" ,
"111111111111110010" , "111111111111111100" , "000000000000000110" , "000000000000001111" , "000000000000011000" , "000000000000100000" , "000000000000100111" , "000000000000101110" , "000000000000110101" , "000000000000111011" ,
"000000000001000001" , "000000000001000110" , "000000000001001011" , "000000000001010000" , "000000000001010100" , "000000000001010111" , "000000000001011011" , "000000000001011110" , "000000000001100000" , "000000000001100010" ,
"000000000001100100" , "000000000001100110" , "000000000001100111" , "000000000001101000" , "000000000001101001" , "000000000001101001" , "000000000001101010" , "000000000001101010" , "000000000001101001" , "000000000001101001" ,
"000000000001101000" , "000000000001101000" , "000000000001100111" , "000000000001100101" , "000000000001100100" , "000000000001100011" , "000000000001100001" , "000000000001011111" , "000000000001011101" , "000000000001011100" ,
"000000000001011010" , "000000000001010111" , "000000000001010101" , "000000000001010011" , "000000000001010001" , "000000000001001110" , "000000000001001100" , "000000000001001010" , "000000000001000111" , "000000000001000101" ,
"000000000001000010" , "000000000001000000" , "000000000000111110" , "000000000000111011" , "000000000000111001" , "000000000000110110" , "000000000000110100" , "000000000000110010" , "000000000000101111" , "000000000000101101" ,
"000000000000101011" , "000000000000101001" , "000000000000100111" , "000000000000100100" , "000000000000100010" , "000000000000100000" , "000000000000011111" , "000000000000011101" , "000000000000011011" , "000000000000011001" ,
"000000000000010111" , "000000000000010110" , "000000000000010100" , "000000000000010011" , "000000000000010001" , "000000000000010000" , "000000000000001111" , "000000000000001101" , "000000000000001100" , "000000000000001011" ,
"000000000000001010" , "000000000000001001" , "000000000000001000" , "000000000000000111" , "000000000000000110" , "000000000000000101" , "000000000000000101" , "000000000000000100" , "000000000000000011" , "000000000000000011" ,
"000000000000000010" , "000000000000000001" , "000000000000000001" , "000000000000000001" , "000000000000000000" , "000000000000000000" , "111111111111111111" , "111111111111111111" , "111111111111111111" , "111111111111111111" ,
"111111111111111111" , "111111111111111110" , "111111111111111110" , "111111111111111110" , "111111111111111110" , "111111111111111110" , "111111111111111110" , "111111111111111110" , "111111111111111110" , "111111111111111110" ,
"111111111111111110" , "111111111111111110" , "111111111111111110" , "111111111111111110" , "111111111111111110" , "111111111111111110" , "111111111111111110" , "111111111111111110" , "111111111111111110" , "111111111111111110" ,
"111111111111111111" , "111111111111111111" , "111111111111111111" , "111111111111111111" , "111111111111111111" , "111111111111111111" , "111111111111111111" , "111111111111111111" , "111111111111111111" , "111111111111111111" ,
"111111111111111111" , "111111111111111111" , "111111111111111111" , "111111111111111111" , "111111111111111111" , "000000000000000000" , "000000000000000000" , "000000000000000000" , "000000000000000000" , "000000000000000000" ,
"000000000000000000" , "000000000000000000" , "000000000000000000" , "000000000000000000" 
);
end a;

