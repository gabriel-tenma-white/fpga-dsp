

library ieee;
library work;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
use work.fft_types.all;

-- delay is 5 cycles

entity windowMultiply1024_64 is
	generic(dataBits, outBits: integer := 18);
	port(clk: in std_logic;
			din: in complex;
			index: in unsigned(10-1 downto 0);
			dout: out complex
			);
end entity;
architecture a of windowMultiply1024_64 is
	constant romDepthOrder: integer := 10;
	constant romDepth: integer := 2**romDepthOrder;
	constant romWidth: integer := 18;
	--ram
	type ram1t is array(0 to romDepth-1) of
		std_logic_vector(romWidth-1 downto 0);
	signal rom: ram1t;
	signal addr1: unsigned(romDepthOrder-1 downto 0);
	signal data0, data1, data2: std_logic_vector(romWidth-1 downto 0);
	signal coeff: signed(romWidth-1 downto 0);

	signal din1, din2, din3: complex;

	-- multiplier
	signal multOutRe, multOutIm: signed(dataBits+romWidth-1 downto 0);
	signal multOut, multOut1: complex;

	attribute keep: string;
	attribute keep of din2: signal is "true";
	attribute keep of data2: signal is "true";
begin
	-- coefficient rom
	addr1 <= index; -- when rising_edge(clk);
	data0 <= rom(to_integer(addr1));
	data1 <= data0 when rising_edge(clk);
	data2 <= data1 when rising_edge(clk);
	coeff <= signed(data2) when rising_edge(clk);

	-- delay data
	din1 <= din when rising_edge(clk);
	din2 <= din1 when rising_edge(clk);
	din3 <= din2 when rising_edge(clk);

	-- multiply
	multOutRe <= coeff * complex_re(din3, dataBits);
	multOutIm <= coeff * complex_im(din3, dataBits);

	multOut <= to_complex(multOutRe(multOutRe'left downto multOutRe'left-outBits+1),
						multOutIm(multOutIm'left downto multOutIm'left-outBits+1));
	multOut1 <= multOut when rising_edge(clk);
	dout <= multOut1 when rising_edge(clk);

	-- rom
	rom <= (

"000000000000000000" , "111111111111100111" , "000000000000000000" , "000000000000110110" , "000000000001000100" , "000000000000010101" , "111111111111011110" , "111111111111010000" , "111111111111100000" , "111111111111100111" ,
"111111111111011110" , "111111111111010111" , "111111111111011001" , "111111111111011001" , "111111111111010010" , "111111111111001100" , "111111111111001010" , "111111111111000111" , "111111111110111111" , "111111111110111000" ,
"111111111110110011" , "111111111110101101" , "111111111110100101" , "111111111110011100" , "111111111110010101" , "111111111110001110" , "111111111110000100" , "111111111101111010" , "111111111101110001" , "111111111101100111" ,
"111111111101011011" , "111111111101001111" , "111111111101000100" , "111111111100111000" , "111111111100101010" , "111111111100011100" , "111111111100001110" , "111111111011111111" , "111111111011101111" , "111111111011011111" ,
"111111111011001111" , "111111111010111101" , "111111111010101011" , "111111111010011000" , "111111111010000101" , "111111111001110001" , "111111111001011100" , "111111111001000110" , "111111111000101111" , "111111111000011001" ,
"111111111000000001" , "111111110111101000" , "111111110111001111" , "111111110110110101" , "111111110110011010" , "111111110101111110" , "111111110101100001" , "111111110101000100" , "111111110100100110" , "111111110100000111" ,
"111111110011101000" , "111111110011000111" , "111111110010100110" , "111111110010000100" , "111111110001100001" , "111111110000111101" , "111111110000011001" , "111111101111110011" , "111111101111001101" , "111111101110100111" ,
"111111101101111111" , "111111101101010111" , "111111101100101110" , "111111101100000100" , "111111101011011001" , "111111101010101110" , "111111101010000010" , "111111101001010101" , "111111101000101000" , "111111100111111010" ,
"111111100111001011" , "111111100110011100" , "111111100101101100" , "111111100100111100" , "111111100100001011" , "111111100011011010" , "111111100010101000" , "111111100001110101" , "111111100001000010" , "111111100000001111" ,
"111111011111011100" , "111111011110101000" , "111111011101110011" , "111111011100111111" , "111111011100001010" , "111111011011010101" , "111111011010100000" , "111111011001101011" , "111111011000110110" , "111111011000000001" ,
"111111010111001100" , "111111010110010111" , "111111010101100001" , "111111010100101101" , "111111010011111000" , "111111010011000100" , "111111010010010000" , "111111010001011100" , "111111010000101001" , "111111001111110111" ,
"111111001111000101" , "111111001110010011" , "111111001101100011" , "111111001100110011" , "111111001100000100" , "111111001011010101" , "111111001010101000" , "111111001001111100" , "111111001001010001" , "111111001000100110" ,
"111111000111111101" , "111111000111010110" , "111111000110101111" , "111111000110001011" , "111111000101100111" , "111111000101000101" , "111111000100100101" , "111111000100000110" , "111111000011101001" , "111111000011001110" ,
"111111000010110101" , "111111000010011110" , "111111000010001001" , "111111000001110110" , "111111000001100101" , "111111000001010110" , "111111000001001010" , "111111000001000000" , "111111000000111000" , "111111000000110011" ,
"111111000000110001" , "111111000000110001" , "111111000000110100" , "111111000000111001" , "111111000001000010" , "111111000001001101" , "111111000001011011" , "111111000001101100" , "111111000010000001" , "111111000010011000" ,
"111111000010110011" , "111111000011010000" , "111111000011110001" , "111111000100010110" , "111111000100111101" , "111111000101101000" , "111111000110010110" , "111111000111001000" , "111111000111111110" , "111111001000110111" ,
"111111001001110011" , "111111001010110011" , "111111001011110111" , "111111001100111110" , "111111001110001001" , "111111001111010111" , "111111010000101001" , "111111010001111111" , "111111010011011001" , "111111010100110110" ,
"111111010110010111" , "111111010111111011" , "111111011001100100" , "111111011011001111" , "111111011100111111" , "111111011110110010" , "111111100000101001" , "111111100010100011" , "111111100100100000" , "111111100110100010" ,
"111111101000100110" , "111111101010101110" , "111111101100111010" , "111111101111001000" , "111111110001011010" , "111111110011101111" , "111111110110000111" , "111111111000100011" , "111111111011000001" , "111111111101100010" ,
"000000000000000101" , "000000000010101100" , "000000000101010101" , "000000001000000001" , "000000001010101111" , "000000001101011111" , "000000010000010001" , "000000010011000110" , "000000010101111100" , "000000011000110101" ,
"000000011011101111" , "000000011110101010" , "000000100001100111" , "000000100100100101" , "000000100111100101" , "000000101010100101" , "000000101101100111" , "000000110000101000" , "000000110011101011" , "000000110110101110" ,
"000000111001110001" , "000000111100110100" , "000000111111110111" , "000001000010111001" , "000001000101111011" , "000001001000111101" , "000001001011111101" , "000001001110111101" , "000001010001111011" , "000001010100111000" ,
"000001010111110011" , "000001011010101100" , "000001011101100011" , "000001100000011000" , "000001100011001011" , "000001100101111011" , "000001101000101000" , "000001101011010010" , "000001101101111000" , "000001110000011100" ,
"000001110010111011" , "000001110101010111" , "000001110111101110" , "000001111010000001" , "000001111100010000" , "000001111110011001" , "000010000000011110" , "000010000010011110" , "000010000100011000" , "000010000110001101" ,
"000010000111111100" , "000010001001100101" , "000010001011001000" , "000010001100100100" , "000010001101111010" , "000010001111001001" , "000010010000010001" , "000010010001010010" , "000010010010001011" , "000010010010111101" ,
"000010010011101000" , "000010010100001010" , "000010010100100101" , "000010010100110111" , "000010010101000001" , "000010010101000010" , "000010010100111010" , "000010010100101010" , "000010010100010001" , "000010010011101111" ,
"000010010011000011" , "000010010010001111" , "000010010001010000" , "000010010000001001" , "000010001110110111" , "000010001101011100" , "000010001011110111" , "000010001010001000" , "000010001000001111" , "000010000110001101" ,
"000010000100000000" , "000010000001101001" , "000001111111000111" , "000001111100011100" , "000001111001100110" , "000001110110100110" , "000001110011011100" , "000001110000001000" , "000001101100101010" , "000001101001000001" ,
"000001100101001111" , "000001100001010010" , "000001011101001011" , "000001011000111011" , "000001010100100000" , "000001001111111100" , "000001001011001110" , "000001000110010111" , "000001000001010110" , "000000111100001100" ,
"000000110110111001" , "000000110001011101" , "000000101011111000" , "000000100110001011" , "000000100000010101" , "000000011010010111" , "000000010100010001" , "000000001110000011" , "000000000111101101" , "000000000001010000" ,
"111111111010101100" , "111111110100000010" , "111111101101010000" , "111111100110011001" , "111111011111011011" , "111111011000011000" , "111111010001010000" , "111111001010000011" , "111111000010110001" , "111110111011011011" ,
"111110110100000001" , "111110101100100011" , "111110100101000010" , "111110011101011110" , "111110010101111000" , "111110001110010000" , "111110000110100110" , "111101111110111100" , "111101110111010000" , "111101101111100100" ,
"111101100111111001" , "111101100000001110" , "111101011000100100" , "111101010000111011" , "111101001001010101" , "111101000001110001" , "111100111010010000" , "111100110010110011" , "111100101011011001" , "111100100100000100" ,
"111100011100110100" , "111100010101101010" , "111100001110100101" , "111100000111100111" , "111100000000110000" , "111011111010000001" , "111011110011011010" , "111011101100111011" , "111011100110100110" , "111011100000011010" ,
"111011011010011001" , "111011010100100010" , "111011001110110110" , "111011001001010111" , "111011000100000100" , "111010111110111101" , "111010111010000100" , "111010110101011001" , "111010110000111101" , "111010101100101111" ,
"111010101000110001" , "111010100101000011" , "111010100001100110" , "111010011110011001" , "111010011011011110" , "111010011000110101" , "111010010110011111" , "111010010100011100" , "111010010010101100" , "111010010001001111" ,
"111010010000001000" , "111010001111010101" , "111010001110110111" , "111010001110101111" , "111010001110111101" , "111010001111100001" , "111010010000011101" , "111010010001101111" , "111010010011011001" , "111010010101011100" ,
"111010010111110110" , "111010011010101001" , "111010011101110110" , "111010100001011011" , "111010100101011010" , "111010101001110011" , "111010101110100110" , "111010110011110100" , "111010111001011100" , "111010111111011111" ,
"111011000101111100" , "111011001100110110" , "111011010100001010" , "111011011011111010" , "111011100100000110" , "111011101100101101" , "111011110101110000" , "111011111111001111" , "111100001001001010" , "111100010011100010" ,
"111100011110010101" , "111100101001100100" , "111100110101001111" , "111101000001010111" , "111101001101111010" , "111101011010111001" , "111101101000010100" , "111101110110001010" , "111110000100011100" , "111110010011001010" ,
"111110100010010010" , "111110110001110110" , "111111000001110100" , "111111010010001101" , "111111100011000000" , "111111110100001101" , "000000000101110100" , "000000010111110100" , "000000101010001101" , "000000111100111111" ,
"000001010000001001" , "000001100011101100" , "000001110111100101" , "000010001011110110" , "000010100000011101" , "000010110101011011" , "000011001010101110" , "000011100000010110" , "000011110110010011" , "000100001100100100" ,
"000100100011001000" , "000100111010000000" , "000101010001001001" , "000101101000100101" , "000110000000010001" , "000110011000001110" , "000110110000011010" , "000111001000110110" , "000111100001100000" , "000111111010011000" ,
"001000010011011100" , "001000101100101101" , "001001000110001001" , "001001011111110000" , "001001111001100001" , "001010010011011011" , "001010101101011101" , "001011000111100111" , "001011100001110111" , "001011111100001110" ,
"001100010110101001" , "001100110001001001" , "001101001011101011" , "001101100110010001" , "001110000000110111" , "001110011011011111" , "001110110110000110" , "001111010000101101" , "001111101011010001" , "010000000101110010" ,
"010000100000010000" , "010000111010101001" , "010001010100111101" , "010001101111001010" , "010010001001001111" , "010010100011001100" , "010010111101000000" , "010011010110101010" , "010011110000001001" , "010100001001011100" ,
"010100100010100011" , "010100111011011011" , "010101010100000101" , "010101101100011111" , "010110000100101001" , "010110011100100010" , "010110110100001001" , "010111001011011100" , "010111100010011100" , "010111111001000111" ,
"011000001111011101" , "011000100101011100" , "011000111011000101" , "011001010000010101" , "011001100101001100" , "011001111001101010" , "011010001101101110" , "011010100001010111" , "011010110100100100" , "011011000111010100" ,
"011011011001100111" , "011011101011011101" , "011011111100110100" , "011100001101101011" , "011100011110000011" , "011100101101111010" , "011100111101010001" , "011101001100000101" , "011101011010011000" , "011101101000000111" ,
"011101110101010011" , "011110000001111100" , "011110001110000000" , "011110011001011111" , "011110100100011010" , "011110101110101110" , "011110111000011101" , "011111000001100101" , "011111001010000111" , "011111010010000001" ,
"011111011001010100" , "011111011111111111" , "011111100110000011" , "011111101011011110" , "011111110000010001" , "011111110100011011" , "011111110111111101" , "011111111010110110" , "011111111101000110" , "011111111110101101" ,
"011111111111101010" , "011111111111111111" , "011111111111101010" , "011111111110101101" , "011111111101000110" , "011111111010110110" , "011111110111111101" , "011111110100011011" , "011111110000010001" , "011111101011011110" ,
"011111100110000011" , "011111011111111111" , "011111011001010100" , "011111010010000001" , "011111001010000111" , "011111000001100101" , "011110111000011101" , "011110101110101110" , "011110100100011010" , "011110011001011111" ,
"011110001110000000" , "011110000001111100" , "011101110101010011" , "011101101000000111" , "011101011010011000" , "011101001100000101" , "011100111101010001" , "011100101101111010" , "011100011110000011" , "011100001101101011" ,
"011011111100110100" , "011011101011011101" , "011011011001100111" , "011011000111010100" , "011010110100100100" , "011010100001010111" , "011010001101101110" , "011001111001101010" , "011001100101001100" , "011001010000010101" ,
"011000111011000101" , "011000100101011100" , "011000001111011101" , "010111111001000111" , "010111100010011100" , "010111001011011100" , "010110110100001001" , "010110011100100010" , "010110000100101001" , "010101101100011111" ,
"010101010100000101" , "010100111011011011" , "010100100010100011" , "010100001001011100" , "010011110000001001" , "010011010110101010" , "010010111101000000" , "010010100011001100" , "010010001001001111" , "010001101111001010" ,
"010001010100111101" , "010000111010101001" , "010000100000010000" , "010000000101110010" , "001111101011010001" , "001111010000101101" , "001110110110000110" , "001110011011011111" , "001110000000110111" , "001101100110010001" ,
"001101001011101011" , "001100110001001001" , "001100010110101001" , "001011111100001110" , "001011100001110111" , "001011000111100111" , "001010101101011101" , "001010010011011011" , "001001111001100001" , "001001011111110000" ,
"001001000110001001" , "001000101100101101" , "001000010011011100" , "000111111010011000" , "000111100001100000" , "000111001000110110" , "000110110000011010" , "000110011000001110" , "000110000000010001" , "000101101000100101" ,
"000101010001001001" , "000100111010000000" , "000100100011001000" , "000100001100100100" , "000011110110010011" , "000011100000010110" , "000011001010101110" , "000010110101011011" , "000010100000011101" , "000010001011110110" ,
"000001110111100101" , "000001100011101100" , "000001010000001001" , "000000111100111111" , "000000101010001101" , "000000010111110100" , "000000000101110100" , "111111110100001101" , "111111100011000000" , "111111010010001101" ,
"111111000001110100" , "111110110001110110" , "111110100010010010" , "111110010011001010" , "111110000100011100" , "111101110110001010" , "111101101000010100" , "111101011010111001" , "111101001101111010" , "111101000001010111" ,
"111100110101001111" , "111100101001100100" , "111100011110010101" , "111100010011100010" , "111100001001001010" , "111011111111001111" , "111011110101110000" , "111011101100101101" , "111011100100000110" , "111011011011111010" ,
"111011010100001010" , "111011001100110110" , "111011000101111100" , "111010111111011111" , "111010111001011100" , "111010110011110100" , "111010101110100110" , "111010101001110011" , "111010100101011010" , "111010100001011011" ,
"111010011101110110" , "111010011010101001" , "111010010111110110" , "111010010101011100" , "111010010011011001" , "111010010001101111" , "111010010000011101" , "111010001111100001" , "111010001110111101" , "111010001110101111" ,
"111010001110110111" , "111010001111010101" , "111010010000001000" , "111010010001001111" , "111010010010101100" , "111010010100011100" , "111010010110011111" , "111010011000110101" , "111010011011011110" , "111010011110011001" ,
"111010100001100110" , "111010100101000011" , "111010101000110001" , "111010101100101111" , "111010110000111101" , "111010110101011001" , "111010111010000100" , "111010111110111101" , "111011000100000100" , "111011001001010111" ,
"111011001110110110" , "111011010100100010" , "111011011010011001" , "111011100000011010" , "111011100110100110" , "111011101100111011" , "111011110011011010" , "111011111010000001" , "111100000000110000" , "111100000111100111" ,
"111100001110100101" , "111100010101101010" , "111100011100110100" , "111100100100000100" , "111100101011011001" , "111100110010110011" , "111100111010010000" , "111101000001110001" , "111101001001010101" , "111101010000111011" ,
"111101011000100100" , "111101100000001110" , "111101100111111001" , "111101101111100100" , "111101110111010000" , "111101111110111100" , "111110000110100110" , "111110001110010000" , "111110010101111000" , "111110011101011110" ,
"111110100101000010" , "111110101100100011" , "111110110100000001" , "111110111011011011" , "111111000010110001" , "111111001010000011" , "111111010001010000" , "111111011000011000" , "111111011111011011" , "111111100110011001" ,
"111111101101010000" , "111111110100000010" , "111111111010101100" , "000000000001010000" , "000000000111101101" , "000000001110000011" , "000000010100010001" , "000000011010010111" , "000000100000010101" , "000000100110001011" ,
"000000101011111000" , "000000110001011101" , "000000110110111001" , "000000111100001100" , "000001000001010110" , "000001000110010111" , "000001001011001110" , "000001001111111100" , "000001010100100000" , "000001011000111011" ,
"000001011101001011" , "000001100001010010" , "000001100101001111" , "000001101001000001" , "000001101100101010" , "000001110000001000" , "000001110011011100" , "000001110110100110" , "000001111001100110" , "000001111100011100" ,
"000001111111000111" , "000010000001101001" , "000010000100000000" , "000010000110001101" , "000010001000001111" , "000010001010001000" , "000010001011110111" , "000010001101011100" , "000010001110110111" , "000010010000001001" ,
"000010010001010000" , "000010010010001111" , "000010010011000011" , "000010010011101111" , "000010010100010001" , "000010010100101010" , "000010010100111010" , "000010010101000010" , "000010010101000001" , "000010010100110111" ,
"000010010100100101" , "000010010100001010" , "000010010011101000" , "000010010010111101" , "000010010010001011" , "000010010001010010" , "000010010000010001" , "000010001111001001" , "000010001101111010" , "000010001100100100" ,
"000010001011001000" , "000010001001100101" , "000010000111111100" , "000010000110001101" , "000010000100011000" , "000010000010011110" , "000010000000011110" , "000001111110011001" , "000001111100010000" , "000001111010000001" ,
"000001110111101110" , "000001110101010111" , "000001110010111011" , "000001110000011100" , "000001101101111000" , "000001101011010010" , "000001101000101000" , "000001100101111011" , "000001100011001011" , "000001100000011000" ,
"000001011101100011" , "000001011010101100" , "000001010111110011" , "000001010100111000" , "000001010001111011" , "000001001110111101" , "000001001011111101" , "000001001000111101" , "000001000101111011" , "000001000010111001" ,
"000000111111110111" , "000000111100110100" , "000000111001110001" , "000000110110101110" , "000000110011101011" , "000000110000101000" , "000000101101100111" , "000000101010100101" , "000000100111100101" , "000000100100100101" ,
"000000100001100111" , "000000011110101010" , "000000011011101111" , "000000011000110101" , "000000010101111100" , "000000010011000110" , "000000010000010001" , "000000001101011111" , "000000001010101111" , "000000001000000001" ,
"000000000101010101" , "000000000010101100" , "000000000000000101" , "111111111101100010" , "111111111011000001" , "111111111000100011" , "111111110110000111" , "111111110011101111" , "111111110001011010" , "111111101111001000" ,
"111111101100111010" , "111111101010101110" , "111111101000100110" , "111111100110100010" , "111111100100100000" , "111111100010100011" , "111111100000101001" , "111111011110110010" , "111111011100111111" , "111111011011001111" ,
"111111011001100100" , "111111010111111011" , "111111010110010111" , "111111010100110110" , "111111010011011001" , "111111010001111111" , "111111010000101001" , "111111001111010111" , "111111001110001001" , "111111001100111110" ,
"111111001011110111" , "111111001010110011" , "111111001001110011" , "111111001000110111" , "111111000111111110" , "111111000111001000" , "111111000110010110" , "111111000101101000" , "111111000100111101" , "111111000100010110" ,
"111111000011110001" , "111111000011010000" , "111111000010110011" , "111111000010011000" , "111111000010000001" , "111111000001101100" , "111111000001011011" , "111111000001001101" , "111111000001000010" , "111111000000111001" ,
"111111000000110100" , "111111000000110001" , "111111000000110001" , "111111000000110011" , "111111000000111000" , "111111000001000000" , "111111000001001010" , "111111000001010110" , "111111000001100101" , "111111000001110110" ,
"111111000010001001" , "111111000010011110" , "111111000010110101" , "111111000011001110" , "111111000011101001" , "111111000100000110" , "111111000100100101" , "111111000101000101" , "111111000101100111" , "111111000110001011" ,
"111111000110101111" , "111111000111010110" , "111111000111111101" , "111111001000100110" , "111111001001010001" , "111111001001111100" , "111111001010101000" , "111111001011010101" , "111111001100000100" , "111111001100110011" ,
"111111001101100011" , "111111001110010011" , "111111001111000101" , "111111001111110111" , "111111010000101001" , "111111010001011100" , "111111010010010000" , "111111010011000100" , "111111010011111000" , "111111010100101101" ,
"111111010101100001" , "111111010110010111" , "111111010111001100" , "111111011000000001" , "111111011000110110" , "111111011001101011" , "111111011010100000" , "111111011011010101" , "111111011100001010" , "111111011100111111" ,
"111111011101110011" , "111111011110101000" , "111111011111011100" , "111111100000001111" , "111111100001000010" , "111111100001110101" , "111111100010101000" , "111111100011011010" , "111111100100001011" , "111111100100111100" ,
"111111100101101100" , "111111100110011100" , "111111100111001011" , "111111100111111010" , "111111101000101000" , "111111101001010101" , "111111101010000010" , "111111101010101110" , "111111101011011001" , "111111101100000100" ,
"111111101100101110" , "111111101101010111" , "111111101101111111" , "111111101110100111" , "111111101111001101" , "111111101111110011" , "111111110000011001" , "111111110000111101" , "111111110001100001" , "111111110010000100" ,
"111111110010100110" , "111111110011000111" , "111111110011101000" , "111111110100000111" , "111111110100100110" , "111111110101000100" , "111111110101100001" , "111111110101111110" , "111111110110011010" , "111111110110110101" ,
"111111110111001111" , "111111110111101000" , "111111111000000001" , "111111111000011001" , "111111111000101111" , "111111111001000110" , "111111111001011100" , "111111111001110001" , "111111111010000101" , "111111111010011000" ,
"111111111010101011" , "111111111010111101" , "111111111011001111" , "111111111011011111" , "111111111011101111" , "111111111011111111" , "111111111100001110" , "111111111100011100" , "111111111100101010" , "111111111100111000" ,
"111111111101000100" , "111111111101001111" , "111111111101011011" , "111111111101100111" , "111111111101110001" , "111111111101111010" , "111111111110000100" , "111111111110001110" , "111111111110010101" , "111111111110011100" ,
"111111111110100101" , "111111111110101101" , "111111111110110011" , "111111111110111000" , "111111111110111111" , "111111111111000111" , "111111111111001010" , "111111111111001100" , "111111111111010010" , "111111111111011001" ,
"111111111111011001" , "111111111111010111" , "111111111111011110" , "111111111111100111" , "111111111111100000" , "111111111111010000" , "111111111111011110" , "000000000000010101" , "000000000001000100" , "000000000000110110" ,
"000000000000000000" , "111111111111100111" , "000000000000000000" , "000000000000010101" 
);
end a;

